module top_module (
clk,
output_1
);

/*
 * We define the type of entries and outputs
 */

input clk;
output [15:0] output_1;


/*
 * Here, we declare some signals need it to pass information between modules
 *
 *
 */

 wire kpn_clk;


/*
 * Here, we instantiate the modules
 *
 *
 */
 
 
 
endmodule